module testbench;

    reg a = 0, b = 0, c = 0, d = 0;

    cadeado cad1(aberto, a, b, c, d);

    always #1 begin
        c <= ~c;
    end

    always #2 begin
        d <= ~d;
    end

initial begin
   $dumpvars;

    a <= 1;
    b <= 1;    

    #500;

   $finish; 
end

endmodule